

module ALU (
    ports
);
    
endmodule
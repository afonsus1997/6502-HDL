

parameter mc_END = 0;
parameter mc_INC_DEC_OP = 1;
parameter mc_INC_DEC = 2; //INC_DEC SRW ACCESS
parameter mc_PC_SRW = 3; //PC GETS registered by SRW bus
parameter mc_PC_AD = 4; //PC GETS can write to AD



module top (
    ports
);
    
endmodule